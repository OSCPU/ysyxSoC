module bitrev (
  input  sck,
  input  ss,
  input  mosi,
  output miso
);
  assign miso = 1'b1;
endmodule
