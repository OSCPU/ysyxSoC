module psram(
  input sck,
  input ce_n,
  inout [3:0] dio
);

  assign dio = 4'bz;

endmodule
